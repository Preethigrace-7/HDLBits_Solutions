module top_module( output one );

// Insert your code here
    int fixme=1;
    assign one = fixme;

endmodule
